library verilog;
use verilog.vl_types.all;
entity DE0_test_vlg_vec_tst is
end DE0_test_vlg_vec_tst;
