LIBRARY ieee;
USE ieee.std_logic_1164.ALL;
USE ieee.std_logic_unsigned.ALL;

ENTITY decoder_5_32 IS
	PORT (
		a : IN STD_LOGIC_VECTOR(4 DOWNTO 0);
		en : IN STD_LOGIC;
		f : OUT STD_LOGIC_VECTOR(31 DOWNTO 0)
	);
END decoder_5_32;

ARCHITECTURE decoder_5_32_a OF decoder_5_32 IS

	SIGNAL p : STD_LOGIC_VECTOR(3 DOWNTO 0);

BEGIN

	p <=
		"1111" WHEN en = '1' ELSE
		"1110" WHEN a(4 DOWNTO 3) = "00" ELSE
		"1101" WHEN a(4 DOWNTO 3) = "01" ELSE
		"1011" WHEN a(4 DOWNTO 3) = "10" ELSE
		"0111";

	f(7 DOWNTO 0) <=
	"11111111" WHEN p(0) = '1' ELSE
	"11111110" WHEN a(2 DOWNTO 0) = o"0" ELSE
	"11111101" WHEN a(2 DOWNTO 0) = o"1" ELSE
	"11111011" WHEN a(2 DOWNTO 0) = o"2" ELSE
	"11110111" WHEN a(2 DOWNTO 0) = o"3" ELSE
	"11101111" WHEN a(2 DOWNTO 0) = o"4" ELSE
	"11011111" WHEN a(2 DOWNTO 0) = o"5" ELSE
	"10111111" WHEN a(2 DOWNTO 0) = o"6" ELSE
	"01111111";

	f(15 DOWNTO 8) <=
	"11111111" WHEN p(1) = '1' ELSE
	"11111110" WHEN a(2 DOWNTO 0) = o"0" ELSE
	"11111101" WHEN a(2 DOWNTO 0) = o"1" ELSE
	"11111011" WHEN a(2 DOWNTO 0) = o"2" ELSE
	"11110111" WHEN a(2 DOWNTO 0) = o"3" ELSE
	"11101111" WHEN a(2 DOWNTO 0) = o"4" ELSE
	"11011111" WHEN a(2 DOWNTO 0) = o"5" ELSE
	"10111111" WHEN a(2 DOWNTO 0) = o"6" ELSE
	"01111111";

	f(23 DOWNTO 16) <=
	"11111111" WHEN p(2) = '1' ELSE
	"11111110" WHEN a(2 DOWNTO 0) = o"0" ELSE
	"11111101" WHEN a(2 DOWNTO 0) = o"1" ELSE
	"11111011" WHEN a(2 DOWNTO 0) = o"2" ELSE
	"11110111" WHEN a(2 DOWNTO 0) = o"3" ELSE
	"11101111" WHEN a(2 DOWNTO 0) = o"4" ELSE
	"11011111" WHEN a(2 DOWNTO 0) = o"5" ELSE
	"10111111" WHEN a(2 DOWNTO 0) = o"6" ELSE
	"01111111";

	f(31 DOWNTO 24) <=
	"11111111" WHEN p(3) = '1' ELSE
	"11111110" WHEN a(2 DOWNTO 0) = o"0" ELSE
	"11111101" WHEN a(2 DOWNTO 0) = o"1" ELSE
	"11111011" WHEN a(2 DOWNTO 0) = o"2" ELSE
	"11110111" WHEN a(2 DOWNTO 0) = o"3" ELSE
	"11101111" WHEN a(2 DOWNTO 0) = o"4" ELSE
	"11011111" WHEN a(2 DOWNTO 0) = o"5" ELSE
	"10111111" WHEN a(2 DOWNTO 0) = o"6" ELSE
	"01111111";

END decoder_5_32_a;