LIBRARY ieee;
USE ieee.std_logic_1164.ALL;
USE ieee.std_logic_unsigned.ALL;

ENTITY decoder_3to8 IS
	PORT (
		A : IN STD_LOGIC;
		B : IN STD_LOGIC;
		C : STD_LOGIC;
		F : OUT STD_LOGIC_VECTOR(7 DOWNTO 0)
	);
END decoder_3to8;
ARCHITECTURE decoder_3to8 OF decoder_3to8 IS
	SIGNAL ABC : STD_LOGIC_VECTOR(2 DOWNTO 0);

BEGIN

	ABC <= A & B & C;
	F <= "00000001" WHEN ABC = o"0" ELSE
		"00000010" WHEN ABC = o"1" ELSE
		"00000100" WHEN ABC = o"2" ELSE
		"00001000" WHEN ABC = o"3" ELSE
		"00010000" WHEN ABC = o"4" ELSE
		"00100000" WHEN ABC = o"5" ELSE
		"01000000" WHEN ABC = o"6" ELSE
		"10000000";

END decoder_3to8;