library verilog;
use verilog.vl_types.all;
entity pwm1_vlg_sample_tst is
    port(
        clk             : in     vl_logic;
        sampler_tx      : out    vl_logic
    );
end pwm1_vlg_sample_tst;
