library verilog;
use verilog.vl_types.all;
entity pwm1_vlg_vec_tst is
end pwm1_vlg_vec_tst;
