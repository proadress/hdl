library verilog;
use verilog.vl_types.all;
entity CPU_ON_DE0_vlg_vec_tst is
end CPU_ON_DE0_vlg_vec_tst;
